*******************************************************************************
* CDL netlist
*
* Library : layout
* Top Cell Name: layout
* View Name: layout
* Netlist created: 13.set.2017
*******************************************************************************

*.SCALE METER
*.GLOBAL 

*******************************************************************************
* Library Name: layout
* Cell Name:    layout
* View Name:    layout
*******************************************************************************

.SUBCKT layout
*.PININFO

.ENDS
